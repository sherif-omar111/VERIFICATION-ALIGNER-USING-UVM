`ifndef CFS_ALGN_TYPES_SV
  `define CFS_ALGN_TYPES_SV

  //Virtual interface
  typedef virtual cfs_algn_if cfs_algn_vif;

`endif