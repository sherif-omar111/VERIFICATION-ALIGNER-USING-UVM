`include "cfs_synch.sv"
`include "cfs_synch_fifo.sv"
`include "cfs_rx_ctrl.sv"
`include "cfs_ctrl.sv"
`include "cfs_tx_ctrl.sv"
`include "cfs_edge_detect.sv"
`include "cfs_regs.sv"
`include "cfs_aligner_core.sv"
`include "cfs_aligner.sv"