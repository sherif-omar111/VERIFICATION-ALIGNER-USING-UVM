`ifndef CFS_ALGN_TEST_DEFINES_SV
  `define CFS_ALGN_TEST_DEFINES_SV

  `ifndef CFS_ALGN_TEST_ALGN_DATA_WIDTH
    `define CFS_ALGN_TEST_ALGN_DATA_WIDTH 32
  `endif

`endif